// How to use:					
// 1. Edit the songs on the Enter Song sheet.					
// 2. Select this whole worksheet, copy it, and paste it into a new file.					
// 3. Save the file as song_rom.v.					
					
module song_rom (					
	input clk,				
	input [8:0] addr,				
	output reg [15:0] dout				
);					
					
	wire [15:0] memory [511:0];				
					
	always @(posedge clk)				
		dout = memory[addr];			
					
	assign memory[	  0	] =	{1'd0, 6'd40, 6'd24, 3'd0};	// Note: 4C
	assign memory[	  1	] =	{1'd0, 6'd44, 6'd24, 3'd0};	// Note: 4E
	assign memory[	  2	] =	{1'd0, 6'd47, 6'd24, 3'd0};	// Note: 4G
	assign memory[	  3	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	  4	] =	{1'd0, 6'd39, 6'd24, 3'd0};	// Note: 4B
	assign memory[	  5	] =	{1'd0, 6'd42, 6'd24, 3'd0};	// Note: 4D
	assign memory[	  6	] =	{1'd0, 6'd47, 6'd24, 3'd0};	// Note: 4G
	assign memory[	  7	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	  8	] =	{1'd0, 6'd37, 6'd24, 3'd0};	// Note: 4A
	assign memory[	  9	] =	{1'd0, 6'd40, 6'd24, 3'd0};	// Note: 4C
	assign memory[	 10	] =	{1'd0, 6'd45, 6'd24, 3'd0};	// Note: 4F
	assign memory[	 11	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	 12	] =	{1'd0, 6'd37, 6'd24, 3'd0};	// Note: 4A
	assign memory[	 13	] =	{1'd0, 6'd42, 6'd24, 3'd0};	// Note: 4D
	assign memory[	 14	] =	{1'd0, 6'd45, 6'd24, 3'd0};	// Note: 4F
	assign memory[	 15	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	 16	] =	{1'd0, 6'd39, 6'd24, 3'd0};	// Note: 4B
	assign memory[	 17	] =	{1'd0, 6'd44, 6'd24, 3'd0};	// Note: 4E
	assign memory[	 18	] =	{1'd0, 6'd48, 6'd24, 3'd0};	// Note: 4G#Ab
	assign memory[	 19	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	 20	] =	{1'd0, 6'd25, 6'd24, 3'd0};	// Note: 3A
	assign memory[	 21	] =	{1'd0, 6'd25, 6'd24, 3'd0};	// Note: 3A
	assign memory[	 22	] =	{1'd0, 6'd25, 6'd24, 3'd0};	// Note: 3A
	assign memory[	 23	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	 24	] =	{1'd0, 6'd27, 6'd24, 3'd0};	// Note: 3B
	assign memory[	 25	] =	{1'd0, 6'd27, 6'd24, 3'd0};	// Note: 3B
	assign memory[	 26	] =	{1'd0, 6'd27, 6'd24, 3'd0};	// Note: 3B
	assign memory[	 27	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	 28	] =	{1'd0, 6'd28, 6'd24, 3'd0};	// Note: 3C
	assign memory[	 29	] =	{1'd0, 6'd28, 6'd24, 3'd0};	// Note: 3C
	assign memory[	 30	] =	{1'd0, 6'd28, 6'd24, 3'd0};	// Note: 3C
	assign memory[	 31	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	 32	] =	{1'd0, 6'd25, 6'd24, 3'd0};	// Note: 3A
	assign memory[	 33	] =	{1'd0, 6'd37, 6'd24, 3'd0};	// Note: 4A
	assign memory[	 34	] =	{1'd0, 6'd49, 6'd24, 3'd0};	// Note: 5A
	assign memory[	 35	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	 36	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 37	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 38	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 39	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 40	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 41	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 42	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 43	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 44	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 45	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 46	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 47	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 48	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 49	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 50	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 51	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 52	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 53	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 54	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 55	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 56	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 57	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 58	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 59	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 60	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 61	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 62	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 63	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 64	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 65	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 66	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 67	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 68	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 69	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 70	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 71	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 72	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 73	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 74	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 75	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 76	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 77	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 78	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 79	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 80	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 81	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 82	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 83	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 84	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 85	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 86	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 87	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 88	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 89	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 90	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 91	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 92	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 93	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 94	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 95	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 96	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 97	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 98	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	 99	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	100	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	101	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	102	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	103	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	104	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	105	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	106	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	107	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	108	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	109	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	110	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	111	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	112	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	113	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	114	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	115	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	116	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	117	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	118	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	119	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	120	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	121	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	122	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	123	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	124	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	125	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	126	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	127	] =	{1'd1, 6'd0, 6'd1, 3'd0};	// Note: rest
	assign memory[	128	] =	{1'd0, 6'd49, 6'd24, 3'd0};	// Note: 5A
	assign memory[	129	] =	{1'd0, 6'd53, 6'd24, 3'd0};	// Note: 5C#Db
	assign memory[	130	] =	{1'd0, 6'd56, 6'd24, 3'd0};	// Note: 5E
	assign memory[	131	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	132	] =	{1'd0, 6'd48, 6'd24, 3'd0};	// Note: 4G#Ab
	assign memory[	133	] =	{1'd0, 6'd39, 6'd24, 3'd0};	// Note: 4B
	assign memory[	134	] =	{1'd0, 6'd54, 6'd24, 3'd0};	// Note: 5D
	assign memory[	135	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	136	] =	{1'd0, 6'd46, 6'd36, 3'd0};	// Note: 4F#Gb
	assign memory[	137	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	138	] =	{1'd0, 6'd53, 6'd24, 3'd0};	// Note: 5C#Db
	assign memory[	139	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	140	] =	{1'd0, 6'd49, 6'd12, 3'd0};	// Note: 5A
	assign memory[	141	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	142	] =	{1'd0, 6'd46, 6'd12, 3'd0};	// Note: 4F#Gb
	assign memory[	143	] =	{1'd0, 6'd53, 6'd12, 3'd0};	// Note: 5C#Db
	assign memory[	144	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	145	] =	{1'd0, 6'd51, 6'd24, 3'd0};	// Note: 5B
	assign memory[	146	] =	{1'd0, 6'd44, 6'd12, 3'd0};	// Note: 4E
	assign memory[	147	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	148	] =	{1'd0, 6'd42, 6'd12, 3'd0};	// Note: 4D
	assign memory[	149	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	150	] =	{1'd0, 6'd41, 6'd12, 3'd0};	// Note: 4C#Db
	assign memory[	151	] =	{1'd0, 6'd45, 6'd12, 3'd0};	// Note: 4F
	assign memory[	152	] =	{1'd0, 6'd53, 6'd12, 3'd0};	// Note: 5C#Db
	assign memory[	153	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	154	] =	{1'd0, 6'd49, 6'd24, 3'd0};	// Note: 5A
	assign memory[	155	] =	{1'd0, 6'd46, 6'd24, 3'd0};	// Note: 4F#Gb
	assign memory[	156	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	157	] =	{1'd0, 6'd46, 6'd24, 3'd0};	// Note: 4F#Gb
	assign memory[	158	] =	{1'd0, 6'd42, 6'd24, 3'd0};	// Note: 4D
	assign memory[	159	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	160	] =	{1'd0, 6'd48, 6'd24, 3'd0};	// Note: 4G#Ab
	assign memory[	161	] =	{1'd0, 6'd45, 6'd24, 3'd0};	// Note: 4F
	assign memory[	162	] =	{1'd0, 6'd41, 6'd24, 3'd0};	// Note: 4C#Db
	assign memory[	163	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	164	] =	{1'd0, 6'd49, 6'd6, 3'd0};	// Note: 5A
	assign memory[	165	] =	{1'd0, 6'd46, 6'd6, 3'd0};	// Note: 4F#Gb
	assign memory[	166	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	167	] =	{1'd0, 6'd48, 6'd6, 3'd0};	// Note: 4G#Ab
	assign memory[	168	] =	{1'd0, 6'd45, 6'd6, 3'd0};	// Note: 4F
	assign memory[	169	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	170	] =	{1'd0, 6'd46, 6'd6, 3'd0};	// Note: 4F#Gb
	assign memory[	171	] =	{1'd0, 6'd41, 6'd6, 3'd0};	// Note: 4C#Db
	assign memory[	172	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	173	] =	{1'd0, 6'd48, 6'd6, 3'd0};	// Note: 4G#Ab
	assign memory[	174	] =	{1'd0, 6'd46, 6'd6, 3'd0};	// Note: 4F#Gb
	assign memory[	175	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	176	] =	{1'd0, 6'd46, 6'd12, 3'd0};	// Note: 4F#Gb
	assign memory[	177	] =	{1'd0, 6'd37, 6'd12, 3'd0};	// Note: 4A
	assign memory[	178	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	179	] =	{1'd0, 6'd48, 6'd12, 3'd0};	// Note: 4G#Ab
	assign memory[	180	] =	{1'd0, 6'd51, 6'd12, 3'd0};	// Note: 5B
	assign memory[	181	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	182	] =	{1'd0, 6'd53, 6'd18, 3'd0};	// Note: 5C#Db
	assign memory[	183	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	184	] =	{1'd0, 6'd46, 6'd12, 3'd0};	// Note: 4F#Gb
	assign memory[	185	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	186	] =	{1'd0, 6'd49, 6'd6, 3'd0};	// Note: 5A
	assign memory[	187	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	188	] =	{1'd0, 6'd54, 6'd6, 3'd0};	// Note: 5D
	assign memory[	189	] =	{1'd0, 6'd51, 6'd6, 3'd0};	// Note: 5B
	assign memory[	190	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	191	] =	{1'd0, 6'd46, 6'd12, 3'd0};	// Note: 4F#Gb
	assign memory[	192	] =	{1'd0, 6'd49, 6'd12, 3'd0};	// Note: 5A
	assign memory[	193	] =	{1'd0, 6'd53, 6'd12, 3'd0};	// Note: 5C#Db
	assign memory[	194	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	195	] =	{1'd0, 6'd46, 6'd12, 3'd0};	// Note: 4F#Gb
	assign memory[	196	] =	{1'd0, 6'd53, 6'd12, 3'd0};	// Note: 5C#Db
	assign memory[	197	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	198	] =	{1'd0, 6'd15, 6'd48, 3'd0};	// Note: 2B
	assign memory[	199	] =	{1'd0, 6'd22, 6'd48, 3'd0};	// Note: 2F#Gb
	assign memory[	200	] =	{1'd0, 6'd51, 6'd6, 3'd0};	// Note: 5B
	assign memory[	201	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	202	] =	{1'd0, 6'd49, 6'd6, 3'd0};	// Note: 5A
	assign memory[	203	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	204	] =	{1'd0, 6'd48, 6'd6, 3'd0};	// Note: 4G#Ab
	assign memory[	205	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	206	] =	{1'd0, 6'd49, 6'd6, 3'd0};	// Note: 5A
	assign memory[	207	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	208	] =	{1'd0, 6'd48, 6'd6, 3'd0};	// Note: 4G#Ab
	assign memory[	209	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	210	] =	{1'd0, 6'd46, 6'd6, 3'd0};	// Note: 4F#Gb
	assign memory[	211	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	212	] =	{1'd0, 6'd44, 6'd6, 3'd0};	// Note: 4E
	assign memory[	213	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	214	] =	{1'd0, 6'd42, 6'd6, 3'd0};	// Note: 4D
	assign memory[	215	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	216	] =	{1'd0, 6'd17, 6'd48, 3'd0};	// Note: 2C#Db
	assign memory[	217	] =	{1'd0, 6'd24, 6'd48, 3'd0};	// Note: 2G#Ab
	assign memory[	218	] =	{1'd0, 6'd41, 6'd6, 3'd0};	// Note: 4C#Db
	assign memory[	219	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	220	] =	{1'd0, 6'd39, 6'd6, 3'd0};	// Note: 4B
	assign memory[	221	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	222	] =	{1'd0, 6'd37, 6'd6, 3'd0};	// Note: 4A
	assign memory[	223	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	224	] =	{1'd0, 6'd36, 6'd6, 3'd0};	// Note: 3G#Ab
	assign memory[	225	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	226	] =	{1'd0, 6'd37, 6'd6, 3'd0};	// Note: 4A
	assign memory[	227	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	228	] =	{1'd0, 6'd39, 6'd6, 3'd0};	// Note: 4B
	assign memory[	229	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	230	] =	{1'd0, 6'd41, 6'd6, 3'd0};	// Note: 4C#Db
	assign memory[	231	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	232	] =	{1'd0, 6'd45, 6'd6, 3'd0};	// Note: 4F
	assign memory[	233	] =	{1'd1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	234	] =	{1'd0, 6'd22, 6'd12, 3'd0};	// Note: 2F#Gb
	assign memory[	235	] =	{1'd0, 6'd34, 6'd12, 3'd0};	// Note: 3F#Gb
	assign memory[	236	] =	{1'd0, 6'd46, 6'd12, 3'd0};	// Note: 4F#Gb
	assign memory[	237	] =	{1'd1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	238	] =	{1'd0, 6'd34, 6'd24, 3'd0};	// Note: 3F#Gb
	assign memory[	239	] =	{1'd0, 6'd41, 6'd24, 3'd0};	// Note: 4C#Db
	assign memory[	240	] =	{1'd0, 6'd49, 6'd24, 3'd0};	// Note: 5A
	assign memory[	241	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	242	] =	{1'd0, 6'd33, 6'd24, 3'd0};	// Note: 3F
	assign memory[	243	] =	{1'd0, 6'd41, 6'd24, 3'd0};	// Note: 4C#Db
	assign memory[	244	] =	{1'd0, 6'd48, 6'd24, 3'd0};	// Note: 4G#Ab
	assign memory[	245	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	246	] =	{1'd0, 6'd30, 6'd24, 3'd0};	// Note: 3D
	assign memory[	247	] =	{1'd0, 6'd37, 6'd24, 3'd0};	// Note: 4A
	assign memory[	248	] =	{1'd0, 6'd46, 6'd24, 3'd0};	// Note: 4F#Gb
	assign memory[	249	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	250	] =	{1'd0, 6'd41, 6'd24, 3'd0};	// Note: 4C#Db
	assign memory[	251	] =	{1'd0, 6'd45, 6'd24, 3'd0};	// Note: 4F
	assign memory[	252	] =	{1'd1, 6'd0, 6'd24, 3'd0};	// Note: rest
	assign memory[	253	] =	{1'd0, 6'd34, 6'd48, 3'd0};	// Note: 3F#Gb
	assign memory[	254	] =	{1'd0, 6'd46, 6'd48, 3'd0};	// Note: 4F#Gb
	assign memory[	255	] =	{1'd1, 6'd0, 6'd48, 3'd0};	// Note: rest
endmodule					
